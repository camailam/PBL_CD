module func21(
	input a,b,c,
	output funcc21
);
not not0(a1,a);
not not1(b1,b);
and and0(funcc21,a1,b1,c);
endmodule 
//verifica se a função da interface 2 é a 2