module func20(
	input a,b,c,
	output funcc20
);
not not0(a1,a);
not not1(b1,b);
and and0(funcc20,a1,b1,c);
endmodule 
//verifica se a função da interface 1 é a 2